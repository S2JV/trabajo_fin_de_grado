** Profile: "SCHEMATIC1-bias"  [ C:\Sebas\02-Facultad\PSpice\02 - Volt�metro\005_etapa_uno_compensado_sim\005_etapa_uno_compensado_sim-pspicefiles\schematic1\bias.sim ] 

** Creating circuit file "bias.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\cds_spb_home\cdssetup\OrCAD_PSpiceTIPSpice_Install\23.1.0\PSpice.ini file:
.lib "C:\Users\sebas\OneDrive - alum.uca.es\B - Spice Models\Transistor\BSS138P.lib" 
.lib "C:\Users\sebas\OneDrive - alum.uca.es\B - Spice Models\Transistor\DMG2302.lib" 
.lib "C:\Users\sebas\OneDrive - alum.uca.es\B - Spice Models\Transistor\2N7000.onsemi.lib" 
.lib "C:\Users\sebas\OneDrive - alum.uca.es\B - Spice Models\Transistor\2N7000.nxp.lib" 
.lib "nom_pspti.lib" 
.lib "nom.lib" 
.inc "C:\Users\sebas\OneDrive - alum.uca.es\04 - Proyectos\01 - [GOAL] TFG\Documentaci�n\include.txt" 

*Analysis directives: 
.TRAN  0 100m 0 0.1m 
.OPTIONS ADVCONV
.OPTIONS FILEMODELSEARCH
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
