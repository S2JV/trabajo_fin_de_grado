** Profile: "SCHEMATIC1-bias"  [ c:\users\sebas\onedrive - alum.uca.es\04 - proyectos\01 - [goal] tfg\01 - dise�os\02 - m�dulo medidor\a - estudios\02 - simulaciones y estudios\01 - resistencia de shunt\03_offset_ai_comp\03_offset_ai_comp-pspicefiles\schematic1\bias.sim ] 

** Creating circuit file "bias.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\cds_spb_home\cdssetup\OrCAD_PSpiceTIPSpice_Install\23.1.0\PSpice.ini file:
.lib "nom_pspti.lib" 
.lib "nom.lib" 

*Analysis directives: 
.OPTIONS ADVCONV
.OPTIONS FILEMODELSEARCH
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
